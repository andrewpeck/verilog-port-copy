module reducer # (
  int    N           = 64,
  int    BRANCH_SIZE = N,
  string OP          = "OR"
) (
  input wire         clk,
  input wire [N-1:0] din,
  output reg         dout
);

  //body
  //
endmodule
